library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


--key schedule
package MY_ARRAY is

	type array28 is array(0 to 16) of STD_LOGIC_VECTOR(0 to 27);
	type array47 is array(0 to 16) of STD_LOGIC_VECTOR(0 to 47);
	type array55 is array(0 to 16) of STD_LOGIC_VECTOR(0 to 55);
	
end MY_ARRAY;
